* ------------------------------------------------------------
* piezo_driver_modes_primary_drive_numeric.cir
* Numeric square drive ACROSS PRIMARY -> transformer -> Lseries -> BVD piezo
* Two runs: MODE=0 (10 ms) and MODE=1 (~100 cycles) with .four
* ------------------------------------------------------------

***** USER PARAMETERS (tune these, not used in PULSE to avoid Mac parsing issues) *****
.param  FDRIVE=108k             ; drive frequency (Hz)
.param  N=3.5                   ; turns ratio Ns/Np
.param  Lp=1m                   ; primary inductance (H)
.param  Ls={Lp*(N**2)}          ; secondary inductance (ideal ratio)
.param  Lseries=120u            ; series inductor on secondary

; Piezo BVD starting params
.param  C0=5n                   ; static (parallel) capacitance
.param  fr=108k                 ; series resonance (Hz)
.param  Qm=80                   ; motional Q
.param  k2=0.12                 ; coupling factor squared

; Soft clamp (~70 Vpp => 35 Vpk)
.param  VCLAMP=35
.param  RCL=500

; Small series resistances for realism/numerical stability
.param  RDRV=0.05               ; series between source and primary
.param  RSEC=0.02               ; tiny R in secondary

***** MODE TRICK (0 = normal, 1 = Fourier) *****
.param MODE=0
.step param MODE list 0 1
.param T0     = {1/FDRIVE}
.param TSTOP  = { if(MODE==0, 10m, 100*T0) }   ; 10 ms vs 100 cycles
.param TW     = {5*T0}                          ; last 5 cycles window

***** DRIVE ACROSS PRIMARY (numeric PULSE, no braces) *****
; ±12 V square at 108 kHz; PW=4.62963us, PER=9.25926us
; Source is between NPDRV and NN (across primary). R in series with primary.
VPRI NPDRV NN PULSE(-12 12 0 10n 10n 4.62963u 9.25926u)
RDRV NP NPDRV 0.05

***** MAGNETICS *****
Lpri NP NN {Lp}
Lsec NS 0  {Ls}
K1   Lpri Lsec 0.998
RSEC_NS NS NS2 {RSEC}
; No NN-to-0 bleed: primary loop is self-contained

***** SECONDARY + MATCHING INDUCTOR + PIEZO *****
Lsec_series NS2 P {Lseries}
XDISC P 0 PIEZO_BVD params: C0={C0} fr={fr} Qm={Qm} k2={k2} Rseries=0.05

; Optional soft clamp (limits V(P) ~ VCLAMP pk)
BI_CLAMP P 0 I = max(0, (V(P)-VCLAMP)/RCL)

***** ANALYSES *****
.options plotwinsize=0 reltol=1e-4 abstol=1e-7
.tran 0 {TSTOP} 0 50n

; Always compute Fourier at FDRIVE (works in both steps)
.four {FDRIVE} V(NS) V(P)

***** SAVE / PROBES *****
.save V(NS) V(NS2) V(P) V(NP) V(NN) V(NPDRV) I(Lpri) I(Lsec) I(Lsec_series)

***** MEASUREMENTS (last 5 cycles of each run) *****
; Transformer secondary (pre-inductor)
.meas TRAN VMAX_SEC   MAX V(NS)             FROM={TSTOP-TW} TO={TSTOP}
.meas TRAN VMIN_SEC   MIN V(NS)             FROM={TSTOP-TW} TO={TSTOP}
.meas TRAN VPP_SEC    PARAM VMAX_SEC - VMIN_SEC
.meas TRAN VRMS_SEC   RMS V(NS)             FROM={TSTOP-TW} TO={TSTOP}

; Piezo terminal (after Lseries)
.meas TRAN VMAX_P     MAX V(P)              FROM={TSTOP-TW} TO={TSTOP}
.meas TRAN VMIN_P     MIN V(P)              FROM={TSTOP-TW} TO={TSTOP}
.meas TRAN VPP_PIEZO  PARAM VMAX_P - VMIN_P
.meas TRAN VRMS_PIEZO RMS V(P)              FROM={TSTOP-TW} TO={TSTOP}
.meas TRAN IRMS_PIEZO RMS I(Lsec_series)    FROM={TSTOP-TW} TO={TSTOP}
.meas TRAN VPK_PIEZO  MAX V(P)              FROM={TSTOP-TW} TO={TSTOP}
.meas TRAN IPK_PIEZO  MAX I(Lsec_series)    FROM={TSTOP-TW} TO={TSTOP}

***** PIEZO SUBCIRCUIT (Butterworth–Van Dyke) *****
* Nodes: P N
* Params: C0, fr, Qm, k2, Rseries(>0 enforced)
.subckt PIEZO_BVD P N params: C0=5n fr=108k Qm=80 k2=0.12 Rleak=200Meg Rseries=0.05
.param w0 = 2*pi*fr
.param Cm = { C0 * k2/(1 - k2) }         ; (or use fa formula if you have fa)
.param Lm = { 1/((w0**2)*Cm) }
.param Rm = { w0*Lm/Qm }

; Parallel static branch (nonzero series R enforced)
Rser P P1 {max(Rseries,1u)}
Csh  P1 N  {C0}
Rle  P  N  {Rleak}

; Motional branch (series Rm-Lm-Cm)
Rm_m  P  M1 {Rm}
Lm_m  M1 M2 {Lm}
Cm_m  M2 N  {Cm}
.ends PIEZO_BVD

***** OPTIONAL DESIGN SWEEPS (uncomment to explore) *****
; .step param N list 3 3.25 3.5 3.75 4
; .step param Lseries list 80u 100u 120u 150u 180u 220u

***** END OF FILE *****
